//////////////////////////////////////////////////////////////////////////////////
// Engineer: 
// Create Date: 2025/01/29 17:34:54
// Module Name: formator
//////////////////////////////////////////////////////////////////////////////////
module formator(

    );



endmodule
